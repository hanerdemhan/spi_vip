interface spi_if (
    input logic clk,
    input logic rst_n
);
    logic mosi;
    logic miso;
    logic sclk;
    logic ss_n;
endinterface
